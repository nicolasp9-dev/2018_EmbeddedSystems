library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all; 
use ieee.std_logic_unsigned.all;

entity LCD_controller is
	port (
	
	Clk      :   IN   std_logic;   
    nReset   :   IN   std_logic; 
	  
	--AVALON slave interface
    AVS_CS       :   IN   std_logic;   
    AVS_Rd       :   IN   std_logic;   
    AVS_Wr       :   IN   std_logic;   
    AVS_RDData   :   OUT  std_logic_vector (31 DOWNTO 0); 
    AVS_WRData   :   IN   std_logic_vector (31 DOWNTO 0); 
    AVS_Adr      :   IN   std_logic_vector (1 DOWNTO 0);
	  
	-- AVALON master inteferace
	AVM_Adr			:OUT		std_logic_vector (31 downto 0 );
	--AVM_ByteEnable	:OUT		std_logic_vector (3 downto 0 );
	--AVM_BurstCount	:OUT		std_logic_vector (2 downto 0 );
	AVM_Rd			:OUT		std_logic;
	AVM_ReadData	:OUT		std_logic_vector (31 downto 0 );
	AVM_WaitRequest	:IN		 	std_logic;
   
	-- LCD output interface
    LCD_ON  	  : OUT 	std_logic  := '1';
	LCD_CS_n 	  : OUT		std_logic  :='1';
	LCD_Reset_n   : OUT		std_logic  :='1';
	LCD_RS 	      : OUT		std_logic  :='1';
	LCD_Wr_n      : OUT		std_logic	:='1';
	LCD_Rd_n      : OUT		std_logic	:='1';
	LCD_data 	  : inOUT	std_logic_vector (15 DOWNTO 0)
		);
		
	end LCD_controller;

	---------------------------------------------------------------------------
architecture rtl of LCD_controller is
	
	
	--declare FIFO component
	--FIFO should be generated by Quartus II
	component fifofifo
	PORT
	(
		clock			: IN STD_LOGIC ;
		data			: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		rdreq			: IN STD_LOGIC ;
		sclr			: IN STD_LOGIC ;
		wrreq			: IN STD_LOGIC ;
		almost_full		: OUT STD_LOGIC ;
		empty			: OUT STD_LOGIC ;
		full			: OUT STD_LOGIC ;
		q				: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		usedw			: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
	end component;
	
	
	
	
	--LCD constant and signals
	constant Nr_line					: integer   := 10;--319;
	constant Nr_column					: integer   := 5;--239;
	constant RW_cycle_default_duration	: integer   := 2;
	
	signal   RW_cycle_duration 			: integer   := 0;
	signal   Line_Counter 				: integer 	:=0;
	signal   Column_Counter 			: integer 	:=0;
	
	
	--state machine
	type LCD_controller_SM is (idle, LCD_start_config, LCD_start_display);
	-- state machine init state
	signal LCD_controller_state : LCD_controller_SM := idle;
	
	--state machine
	type LCD_driver_SM is (LCD_config, LCD_send_CMD_add_register, LCD_send_CMD_to_register, LCD_read_dummy, LCD_read_data, idle,end_of_process, LCD_display_new_picture , LCD_display_next_line, LCD_display_line, LCD_display_pixel_1, LCD_display_pixel_2);
	-- state machine init state
	signal LCD_driver_state : LCD_driver_SM := idle;
	
	--state machine	
	type AVM_SM is (idle, reading, end_of_process);
	--state machine init state
	signal AVM_read_state			: AVM_SM 	:= IDLE;
	
	
	
	--registers
	signal State_register		:		std_logic_vector (31 downto 0);
	signal CMD_address_register	:		std_logic_vector (31 downto 0);
	signal CMD_register			:		std_logic_vector (31 downto 0);
	signal Data_address			:		std_logic_vector (31 downto 0);
	
	--FIFO signals
	signal data_from_FIFO		:		std_logic_vector (31 downto 0);
	signal data_to_FIFO			:		std_logic_vector (31 downto 0);
	signal Rd_FIFO				:		std_logic;
	signal Wr_FIFO				:		std_logic;
	signal empty_FIFO			:		std_logic;
	signal full_FIFO			:		std_logic;
	signal is_not_empty_FIFO	:		std_logic;
	--signal used_space_FIFO		:		std_logic_vector (15 downto 0 );
	signal clear_FIFO			:		std_logic;
	
	-- AVM const
	signal AVM_cnt_read 		:		integer :=0;
	
	
	--flag signals to communicate between process
	signal flag_LCD_config_driver				:		std_logic;
	signal flag_LCD_config_driver_done_reading	:		std_logic;
	signal flag_LCD_config_driver_done_writing 	:		std_logic;
	signal flag_done_displaying					:		std_logic;
	signal flag_start_AVM_read					: 		std_logic;
	signal flag_start_display					: 		std_logic;

	--data signals
	signal LCD_data_read		:		std_logic_vector (7 downto 0); 	
	signal AVM_read_Adr			:		std_logic_vector (31 downto 0);



	---------------------------------------------------------------------------
begin
	
	
	
   fifo_inst: fifofifo
	port map (
		clock			=> clk,
		data			=> data_to_FIFO,
		rdreq			=> Rd_FIFO,
		sclr			=> clear_FIFO,
		wrreq			=> Wr_FIFO,
		almost_full		=> is_not_empty_FIFO,
		empty			=> empty_FIFO,
		full			=> full_FIFO,
		q				=> data_from_FIFO,
		usedw			=> open
	);

   WrReg:            -- Write by Avalon slave access 
   Process(Clk, nReset)   
   Begin   
      if nReset = '0' then  

	  
      end if ; 
   end process WrReg ; 
	
---------------------------------------------------------------------------

   RdReg:            -- Read by Avalon slave access 
   Process(Clk,nreset) 
   Begin
		if  nReset = '0' then  -- init state
		
			AVS_RDData <= (others => '0'); 
			
		elsif rising_edge(clk) then
		  
		  if (AVS_CS = '1') and (AVS_Rd = '1') then 
			 case   AVS_Adr   is   
					when   "00"      =>   AVS_RDData (31 downto 0)  <=  State_register;    
					when   "01"      =>   AVS_RDData (31 downto 0)  <=  CMD_address_register; 
					when   "10"      =>   AVS_RDData (31 downto 0)  <=  CMD_register;
					when   "11"      =>   AVS_RDData (31 downto 0)  <=  Data_address; 			
			   
					when   others   =>    AVS_RDData <= (others => '0'); 
			 end   case;   
		  end if;   
		end if;
   end process RdReg; 

---------------------------------------------------------------------------
   LCD_controller:  -- main FSM of the LCD controller
   Process(Clk, nReset)
   Begin
		if nreset = '0' then
		
			-- init state 
			State_register 			<= (others => '0');
			CMD_address_register 	<= (others => '0');
			CMD_register 			<= (others => '0');
			Data_address 			<= (others => '0');
			
			-- init flag signals
			flag_LCD_config_driver <= '0';
			flag_start_display <= '0';
			
			--init fifo signal			
			clear_FIFO <= '0';
			
		elsif rising_edge(clk) then
		

			if (AVS_CS = '1') and (AVS_Wr = '1') then  -- Write by Avalon slave access 

				case   AVS_Adr    is   
					when   "00"      =>   State_register     	   <=   AVS_WRData (31 downto 0);   
					when   "01"      =>   CMD_address_register     <=   AVS_WRData (31 downto 0); 
					when   "10"      =>   CMD_register     		   <=   AVS_WRData (31 downto 0);
					when   "11"      =>   Data_address    	       <=   AVS_WRData (31 downto 0); 

					when   others   =>   null;   
				end   case; 
				
			else
			
			
			
				case LCD_controller_state is
				
					when idle =>
						
						clear_FIFO <= '0';
									
						if flag_LCD_config_driver = '1' or flag_start_display = '1' then --finalize a process by reseting flags
						
							if (flag_LCD_config_driver_done_reading = '1') then 
							
								flag_LCD_config_driver <= '0';
								State_register(1) <= '0';
								CMD_register (7 downto 0) <= LCD_data_read (7 downto 0 );
								
							elsif (flag_LCD_config_driver_done_writing = '1') then 
							
								flag_LCD_config_driver <= '0';
								State_register(0) <= '0';
								
							elsif (flag_done_displaying = '1') then 
							
								flag_start_display <= '0';
								State_register (2) <= '0';
								
							end if;
						else			--start a new task by assigning flags
							if State_register(0) = '1' then --write cmd
							
								LCD_controller_state <= LCD_start_config;
								
							elsif State_register(1) = '1' then -- read cmd
							
								LCD_controller_state <= LCD_start_config;
							
							elsif State_register(2) = '1' then -- start displaying the image
							
								LCD_controller_state <= LCD_start_display;
								
							end if;
						end if;	
						

						
					when  LCD_start_config =>
						
						flag_LCD_config_driver <= '1';
						
						LCD_controller_state <= idle;

					when LCD_start_display =>
	
						flag_start_display <= '1';
						clear_FIFO <= '1';
						LCD_controller_state <= idle;
						
						
					when others => null;
				end case;
			end if;
		end if;
   end process LCD_controller;
   
   
   LCD_driver: -- LCD_config_read state machine
   Process(Clk, nReset, flag_LCD_config_driver) 
    Begin
		if nReset = '0' then
		
			--init LCD signals
			LCD_data(15 downto 0) 	 <= (others => '0');
			LCD_data_read		    <= (others => '0');
			LCD_ON       			 <= '1';
			LCD_CS_n 	    		 <= '1';
			LCD_Reset_n  			 <= '1';
			LCD_RS 	   				 <= '1';
			LCD_Wr_n        		 <= '1';
			LCD_Rd_n	    		 <= '1';
			
			--init FSM
			LCD_driver_state <= idle;
			
			--init flags
			flag_LCD_config_driver_done_reading <= '0';
			flag_LCD_config_driver_done_writing <= '0';
			
			flag_done_displaying <= '0';
			flag_start_AVM_read <= '0';
			
			--reset FIFO  signals
			Rd_FIFO <= '0';
	  
		elsif rising_edge(clk) then
   
			case LCD_driver_state is
			
				when idle =>
					
					
					
					if flag_LCD_config_driver = '1' then
					
						LCD_driver_state <= LCD_config;	
						
					elsif flag_start_display = '1' then 
					
						LCD_driver_state <= LCD_display_new_picture;
						
					end if;
					
				when end_of_process =>
				
					flag_LCD_config_driver_done_reading <= '0';
					flag_LCD_config_driver_done_writing <= '0';
					flag_done_displaying 				<= '0';
					
					LCD_driver_state <= idle;
					
				when LCD_config =>
				
						LCD_CS_n 	  <= '0';
						LCD_RS 	      <= '0';
						LCD_WR_n      <= '0';
						RW_cycle_duration <= 2*RW_cycle_default_duration;
						
						LCD_driver_state <= LCD_send_CMD_add_register;
						
				when LCD_send_CMD_add_register =>
				
					if RW_cycle_duration > 0 then
					
						LCD_DATA (7 downto 0) <= CMD_address_register (7 downto 0);
						RW_cycle_duration <= RW_cycle_duration - 1;
						
						if RW_cycle_duration = RW_cycle_default_duration then 
							LCD_Wr_n <= '1';
						end if;
						
					else 
						LCD_RS 	      <= '1';
						RW_cycle_duration <= 2*RW_cycle_default_duration;
					
						if State_register(0) = '1' then --write cmd
							LCD_Wr_n	  <= '0';
							
							LCD_driver_state <= LCD_send_CMD_to_register;
							
						elsif State_register(1) = '1' then --read cmnd
							LCD_Rd_n <= '0';
							
							LCD_driver_state <= LCD_read_dummy;
						
						end if;
					end if;
						
						
					when LCD_send_CMD_to_register =>
					
						if RW_cycle_duration > 0 then
						
							LCD_DATA (7 downto 0) <= CMD_register (7 downto 0);
							RW_cycle_duration <= RW_cycle_duration - 1;
							
							if RW_cycle_duration = RW_cycle_default_duration then 
								LCD_Wr_n <= '1';
							end if;
							
						else 
		
						LCD_CS_n 	  <= '1';
						
						flag_LCD_config_driver_done_writing <= '1';
						LCD_driver_state <= end_of_process;
											
						end if;
					
					when LCD_read_dummy =>
							
						if RW_cycle_duration > 0 then
							
							RW_cycle_duration <= RW_cycle_duration - 1;
							
							if RW_cycle_duration = RW_cycle_default_duration then 
								LCD_Rd_n <= '1';
							end if;
							
						else 
							LCD_Rd_n <= '0';
							RW_cycle_duration <= 2*RW_cycle_default_duration;
							LCD_driver_state <= LCD_read_data;	
							
						end if;
						
					when LCD_read_data =>
					
						if RW_cycle_duration > 0 then
							LCD_data_read(7 downto 0) <= LCD_DATA (7 downto 0);
							RW_cycle_duration <= RW_cycle_duration - 1;
							
							if RW_cycle_duration = RW_cycle_default_duration then 
								LCD_Rd_n <= '1';
							end if;
							
						else 
							LCD_CS_n 	  <= '1';
							
							flag_LCD_config_driver_done_reading <= '1';
							LCD_driver_state <= end_of_process;								
						end if;
						
						
					when LCD_display_new_picture =>
					
						LCD_CS_n 	  	<= '0';
						LCD_RS 	      	<= '1';
						Line_Counter	<=	0; -- init number of lines
						
						--ask  AM to access memory and fill FIFO 
						flag_start_AVM_read <= '1';
						
						LCD_driver_state <= LCD_display_next_line;
					
					
					when LCD_display_next_line =>
						
						Column_Counter	<=	0; --init nr of column
						
						if Line_Counter < Nr_line then --display next line on LCD
							Line_Counter <= Line_Counter + 1;
							
							LCD_driver_state <= LCD_display_line;
							
						else --image is completed
						
							flag_done_displaying <= '1';
							LCD_driver_state <= end_of_process;
							
						end if;
						
					when LCD_display_line =>
						
						if Column_counter < Nr_column then
						
							LCD_Wr_n <= '0';
							RW_cycle_duration <= 2*RW_cycle_default_duration;
							
							--get new data from FIFO
							if is_not_empty_FIFO = '1' then 
							
								Rd_FIFO <= '1';
								flag_start_AVM_read <= '0';
								
								LCD_driver_state <= LCD_display_pixel_1;
								
							end if;
							
						else
						
							LCD_driver_state <= LCD_display_next_line; --display next line
							
						end if;

						
					when LCD_display_pixel_1 =>
					
						
						
						if RW_cycle_duration > 0 then
						
							LCD_DATA (15 downto 0) <= data_from_FIFO (15 downto 0);
							
							RW_cycle_duration <= RW_cycle_duration - 1;
							
							Rd_FIFO <= '0';
							
							if RW_cycle_duration = RW_cycle_default_duration then 
							
								LCD_Wr_n <= '1';
								
							end if;
							
						else 
						
							RW_cycle_duration <= 2*RW_cycle_default_duration;
							LCD_Wr_n <= '0';
							Column_counter <= Column_Counter + 1;
							
							LCD_driver_state <= LCD_display_pixel_2;
							
						end if;	
						
					when LCD_display_pixel_2 =>
						
						if RW_cycle_duration > 0 then
						
							LCD_DATA (15 downto 0) <= data_from_FIFO (31 downto 16);
							RW_cycle_duration <= RW_cycle_duration - 1;
							
							if RW_cycle_duration = RW_cycle_default_duration then 
							
								LCD_Wr_n <= '1';
								
							end if;
							
						else 
						
							Column_counter <= Column_Counter + 1;
							LCD_driver_state <= LCD_display_line;
							
						end if;	
						
					when others => null;
			end case;
		end if;
   end process LCD_driver;
   
   Avalon_master_read:            -- Write by Avalon slave access 
   Process(Clk, nReset)   
   Begin   
        if nReset = '0' then  

			--AVM_Adr 			<= (others => '0');
			--AVM_ByteEnable 		<= (others => '0');
			--AVM_BurstCount 		<= (others => '0');
			--AVM_Rd 				<= '0';
			AVM_ReadData 		<= (others => '0');
			AVM_read_Adr		<= (others => '0');
			AVM_cnt_read 	<= 0;
			
			--init FSM
			AVM_read_state <= idle;		
			
			--init FIFO may not be used in final design
			empty_FIFO			<= 'Z';
			full_FIFO			<= 'Z';
			is_not_empty_FIFO	<= 'Z';
			data_to_FIFO		<= (others => 'Z');
			data_from_FIFO		<= (others => 'Z');
			
	    elsif rising_edge(clk) then
		
			case AVM_read_state is
			
				when idle =>
					
					if flag_start_AVM_read = '1' then
					
						AVM_read_state  <= reading;
						AVM_read_Adr	<= Data_address;
						AVM_cnt_read 	<= 0;
						
					end if;
				
				when reading => 
				
					if AVM_WaitRequest /= '1' and full_FIFO /= '1' then 
					
						AVM_read_Adr 		<= AVM_read_Adr + 4;  -- add 4 per word read because master use byte addressing
						AVM_cnt_read 		<= AVM_cnt_read + 1;
						
						if AVM_cnt_read =  Nr_line * Nr_column then  -- 320*240 pixels /2 (as 1 word = 2 pixels)
							
							AVM_read_state <= end_of_process;
							
						end if;
						
					end if;
				
				when end_of_process =>
				
					AVM_read_state <= idle;
					
				when   others   =>   null; 
			end case;
		end if ; 
		
   end process Avalon_master_read ; 
   
   -- read when in reading state and fifo not full
    AVM_Rd <= '1' when AVM_read_state = reading and full_FIFO = '0' else '0';
		

   
   -- write into FIFO if FSM is reading and AVM available and fifo not full
   Wr_FIFO <= '1' when AVM_read_state =  reading and AVM_WaitRequest = '0' and full_FIFO = '0' else '0';
   
	-- this maps the internal address directly to the external port
	AVM_Adr <= AVM_read_Adr;
   
end rtl;