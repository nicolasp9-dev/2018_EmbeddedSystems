-- Author: Nicolas Peslerbe | Embedded system course | UART Programmabe Interface
